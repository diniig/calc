module calc

pub fn add(x int, y int) int {
	println('adding {x} and {y}')
	return x + y
}
